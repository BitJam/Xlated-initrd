   1)  Standard
   2)  checkmd5        Kontrollera live-mediums integritet
   3)  checkfs         Kontrollera LiveUSB ext2/3/4 och persistenta filsystem
   4)  toram           Kopiera det komprimerade filsystemet till RAM
   5)  from=usb        Slutför start från en LiveUSB
   6)  nousb2          Koppla från alla usb-2 enheter vid start
   7)  automount       Montera enheter automatiskt när de pluggas in
   8)  mount=usb       ...och montera alla usb-enheter vid start
   9)  mount=all       ...och montera ALLA usb-enheter vid start
  10)  mount=off       Stäng av all extra montering
  11)  hwclock=ask     Få hjälp av systemet att avgöra klockans inställning
  12)  hwclock=utc     Hårdvaru-klockan använder UTC (Endast Linuxsystem)
  13)  hwclock=local   Hårdvaru-klocka använder lokal tid (Windows system)
  14)  private         Ändra lösenord före start
  15)  nostore         Stäng av LiveUSB-lagringsanvändning
  16)  dostore         Enable LiveUSB-Storage feature
  17)  savestate       Spara en del filer vid omstarter (Endast LiveUSB)
  18)  nosavestate     Spara inte filer vid omstarter (Endast LiveUSB)
