   1)  Standard
   2)  persist_all     Save root in RAM, save home on disk (save root at shutdown)
   3)  persist_root    Save root and home in RAM then saved at shutdown
   4)  persist_static  Save root and home on disk with home separate on disk
   5)  p_static_root   Save root and home on disk together
   6)  persist_home    Bara home-persistens
   7)  frugal_persist  Frugal with root in RAM and home on disk
   8)  frugal_root     Frugal with root and home in RAM then saved at shutdown
   9)  frugal_static   Frugal with root on disk and home separate on disk
  10)  f_static_root   Frugal with root and home on disk together
  11)  frugal_home     Frugal med endast home-persistens
  12)  frugal_only     Bara Frugal, ingen persistens
