   1)  Standard
   2)  checkmd5        Kontrollera live-mediums integritet
   3)  checkfs         Check LiveUSB and persistence ext2/3/4 file systems
   4)  toram           Kopiera det komprimerade filsystemet till RAM
   5)  from=usb        Slutför start från en LiveUSB
   6)  from=hd         Finish booting from a hard drive
   7)  nousb2          Koppla från alla usb-2 enheter vid start
   8)  hwclock=ask     Få hjälp av systemet att avgöra klockans inställning
   9)  hwclock=utc     Hårdvaru-klockan använder UTC (Endast Linuxsystem)
  10)  hwclock=local   Hårdvaru-klocka använder lokal tid (Windows system)
  11)  private         Ändra lösenord före start
  12)  nostore         Disable LiveUSB-Storage feature (LiveUSB only)
  13)  dostore         Enable LiveUSB-Storage feature (LiveUSB only)
  14)  savestate       Spara en del filer vid omstarter (Endast LiveUSB)
  15)  nosavestate     Spara inte filer vid omstarter (Endast LiveUSB)
