   1)  Standard
   2)  automount       Montera enheter automatiskt när de pluggas in
   3)  mount=usb       ...och montera alla usb-enheter vid start
   4)  mount=all       ...och montera ALLA usb-enheter vid start
   5)  mount=off       Disable all extra mounting and automounting
